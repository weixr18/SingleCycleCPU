module Decoder5_32(D , DOUT);
     input wire [4:0] D;
     output wire [31:0] DOUT;

	  assign DOUT =  ({32{(D  == 5'b00000)}} & 32'b00000001) | 
             ({32{(D  == 5'b00001)}} & 32'b00000010) | 
             ({32{(D  == 5'b00010)}} & 32'b00000100) | 
             ({32{(D  == 5'b00011)}} & 32'b00001000) | 
             ({32{(D  == 5'b00100)}} & 32'b00010000) | 
             ({32{(D  == 5'b00101)}} & 32'b00100000) | 
             ({32{(D  == 5'b00110)}} & 32'b01000000) | 
             ({32{(D  == 5'b00111)}} & 32'b10000000) | 
				 
             ({32{(D  == 5'b01000)}} & 32'b00000001_00000000) | 
             ({32{(D  == 5'b01001)}} & 32'b00000010_00000000) | 
             ({32{(D  == 5'b01010)}} & 32'b00000100_00000000) | 
             ({32{(D  == 5'b01011)}} & 32'b00001000_00000000) | 
             ({32{(D  == 5'b01100)}} & 32'b00010000_00000000) | 
             ({32{(D  == 5'b01101)}} & 32'b00100000_00000000) | 
             ({32{(D  == 5'b01110)}} & 32'b01000000_00000000) | 
             ({32{(D  == 5'b01111)}} & 32'b10000000_00000000) | 
              
				 ({32{(D  == 5'b10000)}} & 32'b00000001_00000000_00000000) | 
             ({32{(D  == 5'b10001)}} & 32'b00000010_00000000_00000000) | 
             ({32{(D  == 5'b10010)}} & 32'b00000100_00000000_00000000) | 
             ({32{(D  == 5'b10011)}} & 32'b00001000_00000000_00000000) | 
             ({32{(D  == 5'b10100)}} & 32'b00010000_00000000_00000000) | 
             ({32{(D  == 5'b10101)}} & 32'b00100000_00000000_00000000) | 
             ({32{(D  == 5'b10110)}} & 32'b01000000_00000000_00000000) | 
             ({32{(D  == 5'b10111)}} & 32'b10000000_00000000_00000000) | 
				 
				 ({32{(D  == 5'b11000)}} & 32'b00000001_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11001)}} & 32'b00000010_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11010)}} & 32'b00000100_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11011)}} & 32'b00001000_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11100)}} & 32'b00010000_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11101)}} & 32'b00100000_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11110)}} & 32'b01000000_00000000_00000000_00000000) | 
             ({32{(D  == 5'b11111)}} & 32'b10000000_00000000_00000000_00000000) ;
				 
				 
       
endmodule